module ram();

endmodule
